`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 19.11.2025 02:27:35
// Design Name: 
// Module Name: immediate_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module immediate_top (
    input  logic [31:0] instr,        // Input:Instructions from program memory
    input  logic        imm_sel,      // Input:  0 = Instruction type I, 1 = Instruction type S of control unit
    output logic [31:0] imm32,        // Output for instruction type I and S
    output logic [31:0] imm32_branch  //// Output for instruction type B
);
    logic [11:0] imm12_out;           //  Local variable to store 12-bit immediates - Instructions type I
    logic [12:0] imm13_branch_out;    //  Local variable to store 13-bit immediates - Instructions type B
    //Immediate instruction generator module
    immediate_generator imm1 (
        .instr(instr),                     // Instructions from program memory
        .imm_sel(imm_sel),                 // Multiplexer control from control unit 
        .imm12_out(imm12_out),             // Output of I-type and s-type immediates
        .imm13_branch_out(imm13_branch_out)//Output of B-type immediates
    );
 
 // Sign-extension module for I-type and S-type instructions
    extend_sign #(.WIDTH_IN(12), .WIDTH_OUT(32)) extend_i_s (
        .imm_in(imm12_out),       // I-type and S-type immediates generated by the immediate generator module  
        .imm_out(imm32)           //output for  ALU
    );
 // Sign-extension module for B-type instructions
   extend_sign #(.WIDTH_IN(13), .WIDTH_OUT(32)) extend_branch (
        .imm_in(imm13_branch_out),       // B-type immediates generated by the immediate generator module  
        .imm_out(imm32_branch)           //output for  PROGRAM COUNTER
    );

endmodule

