`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/22/2025 02:26:58 AM
// Design Name: 
// Module Name: program_counter
// Project Name: 
//////////////////////////////////////////////////////////////////////////////////

module program_counter(
    input logic clk,
    input logic arst_n,
    input logic pc_write,
    input logic zero,
    input logic [1:0] pc_sel,
    input logic [31:0] pc_imm_in,
    output logic [31:0] pc
);

`include "defines.svh"

    
    //Secuential logic 
    always_ff @(posedge clk, negedge arst_n) begin
        if (!arst_n) begin
            pc <= 32'h0000_0000;
        end else if (pc_write) begin
            unique case (pc_sel)
                PC_4: begin 
                    pc <= pc + 4;        
                end
                PC_BRANCH: begin
                    if (zero) begin  //if branch taken
                        pc <= pc + pc_imm_in; 
                    end else begin 
                        pc <= pc + 4;
                    end
                end
                PC_JAL: begin
                    pc <= pc + pc_imm_in; 
                end  
                default: begin 
                    pc <= pc;
                end    
            endcase
        end 
    end    
endmodule



