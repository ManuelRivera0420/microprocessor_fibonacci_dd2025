module mux #(parameter N = 8) (

	);
	endmodule
