 module microprocessor_tb ();

 endmodule
