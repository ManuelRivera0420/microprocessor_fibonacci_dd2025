module microprocessor (
	
);

endmodule
